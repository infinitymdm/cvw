module fdivsqrtuslc4 (
	Dmsbs,
	Smsbs,
	WSmsbs,
	WCmsbs,
	Sqrt,
	j0,
	j1,
	udigit
);
	reg _sv2v_0;
	input wire [2:0] Dmsbs;
	input wire [4:0] Smsbs;
	input wire [7:0] WSmsbs;
	input wire [7:0] WCmsbs;
	input wire Sqrt;
	input wire j0;
	input wire j1;
	output wire [3:0] udigit;
	wire [7:0] PreWmsbs;
	wire [6:0] Wmsbs;
	reg [2:0] A;
	assign PreWmsbs = WCmsbs + WSmsbs;
	assign Wmsbs = PreWmsbs[7:1];
	reg [3:0] USel4;
	always @(*) begin : sv2v_autoblock_1
		case ({A, Wmsbs})
			10'd0: USel4 = 4'b0000;
			10'd1: USel4 = 4'b0000;
			10'd2: USel4 = 4'b0000;
			10'd3: USel4 = 4'b0000;
			10'd4: USel4 = 4'b0100;
			10'd5: USel4 = 4'b0100;
			10'd6: USel4 = 4'b0100;
			10'd7: USel4 = 4'b0100;
			10'd8: USel4 = 4'b0100;
			10'd9: USel4 = 4'b0100;
			10'd10: USel4 = 4'b0100;
			10'd11: USel4 = 4'b0100;
			10'd12: USel4 = 4'b1000;
			10'd13: USel4 = 4'b1000;
			10'd14: USel4 = 4'b1000;
			10'd15: USel4 = 4'b1000;
			10'd16: USel4 = 4'b1000;
			10'd17: USel4 = 4'b1000;
			10'd18: USel4 = 4'b1000;
			10'd19: USel4 = 4'b1000;
			10'd20: USel4 = 4'b1000;
			10'd21: USel4 = 4'b1000;
			10'd22: USel4 = 4'b1000;
			10'd23: USel4 = 4'b1000;
			10'd24: USel4 = 4'b1000;
			10'd25: USel4 = 4'b1000;
			10'd26: USel4 = 4'b1000;
			10'd27: USel4 = 4'b1000;
			10'd28: USel4 = 4'b1000;
			10'd29: USel4 = 4'b1000;
			10'd30: USel4 = 4'b1000;
			10'd31: USel4 = 4'b1000;
			10'd32: USel4 = 4'b1000;
			10'd33: USel4 = 4'b1000;
			10'd34: USel4 = 4'b1000;
			10'd35: USel4 = 4'b1000;
			10'd36: USel4 = 4'b1000;
			10'd37: USel4 = 4'b1000;
			10'd38: USel4 = 4'b1000;
			10'd39: USel4 = 4'b1000;
			10'd40: USel4 = 4'b1000;
			10'd41: USel4 = 4'b1000;
			10'd42: USel4 = 4'b1000;
			10'd43: USel4 = 4'b1000;
			10'd44: USel4 = 4'b1000;
			10'd45: USel4 = 4'b1000;
			10'd46: USel4 = 4'b1000;
			10'd47: USel4 = 4'b1000;
			10'd48: USel4 = 4'b1000;
			10'd49: USel4 = 4'b1000;
			10'd50: USel4 = 4'b1000;
			10'd51: USel4 = 4'b1000;
			10'd52: USel4 = 4'b1000;
			10'd53: USel4 = 4'b1000;
			10'd54: USel4 = 4'b1000;
			10'd55: USel4 = 4'b1000;
			10'd56: USel4 = 4'b1000;
			10'd57: USel4 = 4'b1000;
			10'd58: USel4 = 4'b1000;
			10'd59: USel4 = 4'b1000;
			10'd60: USel4 = 4'b1000;
			10'd61: USel4 = 4'b1000;
			10'd62: USel4 = 4'b1000;
			10'd63: USel4 = 4'b1000;
			10'd64: USel4 = 4'b0001;
			10'd65: USel4 = 4'b0001;
			10'd66: USel4 = 4'b0001;
			10'd67: USel4 = 4'b0001;
			10'd68: USel4 = 4'b0001;
			10'd69: USel4 = 4'b0001;
			10'd70: USel4 = 4'b0001;
			10'd71: USel4 = 4'b0001;
			10'd72: USel4 = 4'b0001;
			10'd73: USel4 = 4'b0001;
			10'd74: USel4 = 4'b0001;
			10'd75: USel4 = 4'b0001;
			10'd76: USel4 = 4'b0001;
			10'd77: USel4 = 4'b0001;
			10'd78: USel4 = 4'b0001;
			10'd79: USel4 = 4'b0001;
			10'd80: USel4 = 4'b0001;
			10'd81: USel4 = 4'b0001;
			10'd82: USel4 = 4'b0001;
			10'd83: USel4 = 4'b0001;
			10'd84: USel4 = 4'b0001;
			10'd85: USel4 = 4'b0001;
			10'd86: USel4 = 4'b0001;
			10'd87: USel4 = 4'b0001;
			10'd88: USel4 = 4'b0001;
			10'd89: USel4 = 4'b0001;
			10'd90: USel4 = 4'b0001;
			10'd91: USel4 = 4'b0001;
			10'd92: USel4 = 4'b0001;
			10'd93: USel4 = 4'b0001;
			10'd94: USel4 = 4'b0001;
			10'd95: USel4 = 4'b0001;
			10'd96: USel4 = 4'b0001;
			10'd97: USel4 = 4'b0001;
			10'd98: USel4 = 4'b0001;
			10'd99: USel4 = 4'b0001;
			10'd100: USel4 = 4'b0001;
			10'd101: USel4 = 4'b0001;
			10'd102: USel4 = 4'b0001;
			10'd103: USel4 = 4'b0001;
			10'd104: USel4 = 4'b0001;
			10'd105: USel4 = 4'b0001;
			10'd106: USel4 = 4'b0001;
			10'd107: USel4 = 4'b0001;
			10'd108: USel4 = 4'b0001;
			10'd109: USel4 = 4'b0001;
			10'd110: USel4 = 4'b0001;
			10'd111: USel4 = 4'b0001;
			10'd112: USel4 = 4'b0001;
			10'd113: USel4 = 4'b0001;
			10'd114: USel4 = 4'b0001;
			10'd115: USel4 = 4'b0010;
			10'd116: USel4 = 4'b0010;
			10'd117: USel4 = 4'b0010;
			10'd118: USel4 = 4'b0010;
			10'd119: USel4 = 4'b0010;
			10'd120: USel4 = 4'b0010;
			10'd121: USel4 = 4'b0010;
			10'd122: USel4 = 4'b0010;
			10'd123: USel4 = 4'b0010;
			10'd124: USel4 = 4'b0000;
			10'd125: USel4 = 4'b0000;
			10'd126: USel4 = 4'b0000;
			10'd127: USel4 = 4'b0000;
			10'd128: USel4 = 4'b0000;
			10'd129: USel4 = 4'b0000;
			10'd130: USel4 = 4'b0000;
			10'd131: USel4 = 4'b0000;
			10'd132: USel4 = 4'b0100;
			10'd133: USel4 = 4'b0100;
			10'd134: USel4 = 4'b0100;
			10'd135: USel4 = 4'b0100;
			10'd136: USel4 = 4'b0100;
			10'd137: USel4 = 4'b0100;
			10'd138: USel4 = 4'b0100;
			10'd139: USel4 = 4'b0100;
			10'd140: USel4 = 4'b0100;
			10'd141: USel4 = 4'b0100;
			10'd142: USel4 = 4'b1000;
			10'd143: USel4 = 4'b1000;
			10'd144: USel4 = 4'b1000;
			10'd145: USel4 = 4'b1000;
			10'd146: USel4 = 4'b1000;
			10'd147: USel4 = 4'b1000;
			10'd148: USel4 = 4'b1000;
			10'd149: USel4 = 4'b1000;
			10'd150: USel4 = 4'b1000;
			10'd151: USel4 = 4'b1000;
			10'd152: USel4 = 4'b1000;
			10'd153: USel4 = 4'b1000;
			10'd154: USel4 = 4'b1000;
			10'd155: USel4 = 4'b1000;
			10'd156: USel4 = 4'b1000;
			10'd157: USel4 = 4'b1000;
			10'd158: USel4 = 4'b1000;
			10'd159: USel4 = 4'b1000;
			10'd160: USel4 = 4'b1000;
			10'd161: USel4 = 4'b1000;
			10'd162: USel4 = 4'b1000;
			10'd163: USel4 = 4'b1000;
			10'd164: USel4 = 4'b1000;
			10'd165: USel4 = 4'b1000;
			10'd166: USel4 = 4'b1000;
			10'd167: USel4 = 4'b1000;
			10'd168: USel4 = 4'b1000;
			10'd169: USel4 = 4'b1000;
			10'd170: USel4 = 4'b1000;
			10'd171: USel4 = 4'b1000;
			10'd172: USel4 = 4'b1000;
			10'd173: USel4 = 4'b1000;
			10'd174: USel4 = 4'b1000;
			10'd175: USel4 = 4'b1000;
			10'd176: USel4 = 4'b1000;
			10'd177: USel4 = 4'b1000;
			10'd178: USel4 = 4'b1000;
			10'd179: USel4 = 4'b1000;
			10'd180: USel4 = 4'b1000;
			10'd181: USel4 = 4'b1000;
			10'd182: USel4 = 4'b1000;
			10'd183: USel4 = 4'b1000;
			10'd184: USel4 = 4'b1000;
			10'd185: USel4 = 4'b1000;
			10'd186: USel4 = 4'b1000;
			10'd187: USel4 = 4'b1000;
			10'd188: USel4 = 4'b1000;
			10'd189: USel4 = 4'b1000;
			10'd190: USel4 = 4'b1000;
			10'd191: USel4 = 4'b1000;
			10'd192: USel4 = 4'b0001;
			10'd193: USel4 = 4'b0001;
			10'd194: USel4 = 4'b0001;
			10'd195: USel4 = 4'b0001;
			10'd196: USel4 = 4'b0001;
			10'd197: USel4 = 4'b0001;
			10'd198: USel4 = 4'b0001;
			10'd199: USel4 = 4'b0001;
			10'd200: USel4 = 4'b0001;
			10'd201: USel4 = 4'b0001;
			10'd202: USel4 = 4'b0001;
			10'd203: USel4 = 4'b0001;
			10'd204: USel4 = 4'b0001;
			10'd205: USel4 = 4'b0001;
			10'd206: USel4 = 4'b0001;
			10'd207: USel4 = 4'b0001;
			10'd208: USel4 = 4'b0001;
			10'd209: USel4 = 4'b0001;
			10'd210: USel4 = 4'b0001;
			10'd211: USel4 = 4'b0001;
			10'd212: USel4 = 4'b0001;
			10'd213: USel4 = 4'b0001;
			10'd214: USel4 = 4'b0001;
			10'd215: USel4 = 4'b0001;
			10'd216: USel4 = 4'b0001;
			10'd217: USel4 = 4'b0001;
			10'd218: USel4 = 4'b0001;
			10'd219: USel4 = 4'b0001;
			10'd220: USel4 = 4'b0001;
			10'd221: USel4 = 4'b0001;
			10'd222: USel4 = 4'b0001;
			10'd223: USel4 = 4'b0001;
			10'd224: USel4 = 4'b0001;
			10'd225: USel4 = 4'b0001;
			10'd226: USel4 = 4'b0001;
			10'd227: USel4 = 4'b0001;
			10'd228: USel4 = 4'b0001;
			10'd229: USel4 = 4'b0001;
			10'd230: USel4 = 4'b0001;
			10'd231: USel4 = 4'b0001;
			10'd232: USel4 = 4'b0001;
			10'd233: USel4 = 4'b0001;
			10'd234: USel4 = 4'b0001;
			10'd235: USel4 = 4'b0001;
			10'd236: USel4 = 4'b0001;
			10'd237: USel4 = 4'b0001;
			10'd238: USel4 = 4'b0001;
			10'd239: USel4 = 4'b0001;
			10'd240: USel4 = 4'b0001;
			10'd241: USel4 = 4'b0001;
			10'd242: USel4 = 4'b0010;
			10'd243: USel4 = 4'b0010;
			10'd244: USel4 = 4'b0010;
			10'd245: USel4 = 4'b0010;
			10'd246: USel4 = 4'b0010;
			10'd247: USel4 = 4'b0010;
			10'd248: USel4 = 4'b0010;
			10'd249: USel4 = 4'b0010;
			10'd250: USel4 = 4'b0010;
			10'd251: USel4 = 4'b0010;
			10'd252: USel4 = 4'b0000;
			10'd253: USel4 = 4'b0000;
			10'd254: USel4 = 4'b0000;
			10'd255: USel4 = 4'b0000;
			10'd256: USel4 = 4'b0000;
			10'd257: USel4 = 4'b0000;
			10'd258: USel4 = 4'b0000;
			10'd259: USel4 = 4'b0000;
			10'd260: USel4 = 4'b0100;
			10'd261: USel4 = 4'b0100;
			10'd262: USel4 = 4'b0100;
			10'd263: USel4 = 4'b0100;
			10'd264: USel4 = 4'b0100;
			10'd265: USel4 = 4'b0100;
			10'd266: USel4 = 4'b0100;
			10'd267: USel4 = 4'b0100;
			10'd268: USel4 = 4'b0100;
			10'd269: USel4 = 4'b0100;
			10'd270: USel4 = 4'b0100;
			10'd271: USel4 = 4'b0100;
			10'd272: USel4 = 4'b1000;
			10'd273: USel4 = 4'b1000;
			10'd274: USel4 = 4'b1000;
			10'd275: USel4 = 4'b1000;
			10'd276: USel4 = 4'b1000;
			10'd277: USel4 = 4'b1000;
			10'd278: USel4 = 4'b1000;
			10'd279: USel4 = 4'b1000;
			10'd280: USel4 = 4'b1000;
			10'd281: USel4 = 4'b1000;
			10'd282: USel4 = 4'b1000;
			10'd283: USel4 = 4'b1000;
			10'd284: USel4 = 4'b1000;
			10'd285: USel4 = 4'b1000;
			10'd286: USel4 = 4'b1000;
			10'd287: USel4 = 4'b1000;
			10'd288: USel4 = 4'b1000;
			10'd289: USel4 = 4'b1000;
			10'd290: USel4 = 4'b1000;
			10'd291: USel4 = 4'b1000;
			10'd292: USel4 = 4'b1000;
			10'd293: USel4 = 4'b1000;
			10'd294: USel4 = 4'b1000;
			10'd295: USel4 = 4'b1000;
			10'd296: USel4 = 4'b1000;
			10'd297: USel4 = 4'b1000;
			10'd298: USel4 = 4'b1000;
			10'd299: USel4 = 4'b1000;
			10'd300: USel4 = 4'b1000;
			10'd301: USel4 = 4'b1000;
			10'd302: USel4 = 4'b1000;
			10'd303: USel4 = 4'b1000;
			10'd304: USel4 = 4'b1000;
			10'd305: USel4 = 4'b1000;
			10'd306: USel4 = 4'b1000;
			10'd307: USel4 = 4'b1000;
			10'd308: USel4 = 4'b1000;
			10'd309: USel4 = 4'b1000;
			10'd310: USel4 = 4'b1000;
			10'd311: USel4 = 4'b1000;
			10'd312: USel4 = 4'b1000;
			10'd313: USel4 = 4'b1000;
			10'd314: USel4 = 4'b1000;
			10'd315: USel4 = 4'b1000;
			10'd316: USel4 = 4'b1000;
			10'd317: USel4 = 4'b1000;
			10'd318: USel4 = 4'b1000;
			10'd319: USel4 = 4'b1000;
			10'd320: USel4 = 4'b0001;
			10'd321: USel4 = 4'b0001;
			10'd322: USel4 = 4'b0001;
			10'd323: USel4 = 4'b0001;
			10'd324: USel4 = 4'b0001;
			10'd325: USel4 = 4'b0001;
			10'd326: USel4 = 4'b0001;
			10'd327: USel4 = 4'b0001;
			10'd328: USel4 = 4'b0001;
			10'd329: USel4 = 4'b0001;
			10'd330: USel4 = 4'b0001;
			10'd331: USel4 = 4'b0001;
			10'd332: USel4 = 4'b0001;
			10'd333: USel4 = 4'b0001;
			10'd334: USel4 = 4'b0001;
			10'd335: USel4 = 4'b0001;
			10'd336: USel4 = 4'b0001;
			10'd337: USel4 = 4'b0001;
			10'd338: USel4 = 4'b0001;
			10'd339: USel4 = 4'b0001;
			10'd340: USel4 = 4'b0001;
			10'd341: USel4 = 4'b0001;
			10'd342: USel4 = 4'b0001;
			10'd343: USel4 = 4'b0001;
			10'd344: USel4 = 4'b0001;
			10'd345: USel4 = 4'b0001;
			10'd346: USel4 = 4'b0001;
			10'd347: USel4 = 4'b0001;
			10'd348: USel4 = 4'b0001;
			10'd349: USel4 = 4'b0001;
			10'd350: USel4 = 4'b0001;
			10'd351: USel4 = 4'b0001;
			10'd352: USel4 = 4'b0001;
			10'd353: USel4 = 4'b0001;
			10'd354: USel4 = 4'b0001;
			10'd355: USel4 = 4'b0001;
			10'd356: USel4 = 4'b0001;
			10'd357: USel4 = 4'b0001;
			10'd358: USel4 = 4'b0001;
			10'd359: USel4 = 4'b0001;
			10'd360: USel4 = 4'b0001;
			10'd361: USel4 = 4'b0001;
			10'd362: USel4 = 4'b0001;
			10'd363: USel4 = 4'b0001;
			10'd364: USel4 = 4'b0001;
			10'd365: USel4 = 4'b0001;
			10'd366: USel4 = 4'b0001;
			10'd367: USel4 = 4'b0001;
			10'd368: USel4 = 4'b0010;
			10'd369: USel4 = 4'b0010;
			10'd370: USel4 = 4'b0010;
			10'd371: USel4 = 4'b0010;
			10'd372: USel4 = 4'b0010;
			10'd373: USel4 = 4'b0010;
			10'd374: USel4 = 4'b0010;
			10'd375: USel4 = 4'b0010;
			10'd376: USel4 = 4'b0010;
			10'd377: USel4 = 4'b0010;
			10'd378: USel4 = 4'b0000;
			10'd379: USel4 = 4'b0000;
			10'd380: USel4 = 4'b0000;
			10'd381: USel4 = 4'b0000;
			10'd382: USel4 = 4'b0000;
			10'd383: USel4 = 4'b0000;
			10'd384: USel4 = 4'b0000;
			10'd385: USel4 = 4'b0000;
			10'd386: USel4 = 4'b0000;
			10'd387: USel4 = 4'b0000;
			10'd388: USel4 = 4'b0100;
			10'd389: USel4 = 4'b0100;
			10'd390: USel4 = 4'b0100;
			10'd391: USel4 = 4'b0100;
			10'd392: USel4 = 4'b0100;
			10'd393: USel4 = 4'b0100;
			10'd394: USel4 = 4'b0100;
			10'd395: USel4 = 4'b0100;
			10'd396: USel4 = 4'b0100;
			10'd397: USel4 = 4'b0100;
			10'd398: USel4 = 4'b0100;
			10'd399: USel4 = 4'b0100;
			10'd400: USel4 = 4'b1000;
			10'd401: USel4 = 4'b1000;
			10'd402: USel4 = 4'b1000;
			10'd403: USel4 = 4'b1000;
			10'd404: USel4 = 4'b1000;
			10'd405: USel4 = 4'b1000;
			10'd406: USel4 = 4'b1000;
			10'd407: USel4 = 4'b1000;
			10'd408: USel4 = 4'b1000;
			10'd409: USel4 = 4'b1000;
			10'd410: USel4 = 4'b1000;
			10'd411: USel4 = 4'b1000;
			10'd412: USel4 = 4'b1000;
			10'd413: USel4 = 4'b1000;
			10'd414: USel4 = 4'b1000;
			10'd415: USel4 = 4'b1000;
			10'd416: USel4 = 4'b1000;
			10'd417: USel4 = 4'b1000;
			10'd418: USel4 = 4'b1000;
			10'd419: USel4 = 4'b1000;
			10'd420: USel4 = 4'b1000;
			10'd421: USel4 = 4'b1000;
			10'd422: USel4 = 4'b1000;
			10'd423: USel4 = 4'b1000;
			10'd424: USel4 = 4'b1000;
			10'd425: USel4 = 4'b1000;
			10'd426: USel4 = 4'b1000;
			10'd427: USel4 = 4'b1000;
			10'd428: USel4 = 4'b1000;
			10'd429: USel4 = 4'b1000;
			10'd430: USel4 = 4'b1000;
			10'd431: USel4 = 4'b1000;
			10'd432: USel4 = 4'b1000;
			10'd433: USel4 = 4'b1000;
			10'd434: USel4 = 4'b1000;
			10'd435: USel4 = 4'b1000;
			10'd436: USel4 = 4'b1000;
			10'd437: USel4 = 4'b1000;
			10'd438: USel4 = 4'b1000;
			10'd439: USel4 = 4'b1000;
			10'd440: USel4 = 4'b1000;
			10'd441: USel4 = 4'b1000;
			10'd442: USel4 = 4'b1000;
			10'd443: USel4 = 4'b1000;
			10'd444: USel4 = 4'b1000;
			10'd445: USel4 = 4'b1000;
			10'd446: USel4 = 4'b1000;
			10'd447: USel4 = 4'b1000;
			10'd448: USel4 = 4'b0001;
			10'd449: USel4 = 4'b0001;
			10'd450: USel4 = 4'b0001;
			10'd451: USel4 = 4'b0001;
			10'd452: USel4 = 4'b0001;
			10'd453: USel4 = 4'b0001;
			10'd454: USel4 = 4'b0001;
			10'd455: USel4 = 4'b0001;
			10'd456: USel4 = 4'b0001;
			10'd457: USel4 = 4'b0001;
			10'd458: USel4 = 4'b0001;
			10'd459: USel4 = 4'b0001;
			10'd460: USel4 = 4'b0001;
			10'd461: USel4 = 4'b0001;
			10'd462: USel4 = 4'b0001;
			10'd463: USel4 = 4'b0001;
			10'd464: USel4 = 4'b0001;
			10'd465: USel4 = 4'b0001;
			10'd466: USel4 = 4'b0001;
			10'd467: USel4 = 4'b0001;
			10'd468: USel4 = 4'b0001;
			10'd469: USel4 = 4'b0001;
			10'd470: USel4 = 4'b0001;
			10'd471: USel4 = 4'b0001;
			10'd472: USel4 = 4'b0001;
			10'd473: USel4 = 4'b0001;
			10'd474: USel4 = 4'b0001;
			10'd475: USel4 = 4'b0001;
			10'd476: USel4 = 4'b0001;
			10'd477: USel4 = 4'b0001;
			10'd478: USel4 = 4'b0001;
			10'd479: USel4 = 4'b0001;
			10'd480: USel4 = 4'b0001;
			10'd481: USel4 = 4'b0001;
			10'd482: USel4 = 4'b0001;
			10'd483: USel4 = 4'b0001;
			10'd484: USel4 = 4'b0001;
			10'd485: USel4 = 4'b0001;
			10'd486: USel4 = 4'b0001;
			10'd487: USel4 = 4'b0001;
			10'd488: USel4 = 4'b0001;
			10'd489: USel4 = 4'b0001;
			10'd490: USel4 = 4'b0001;
			10'd491: USel4 = 4'b0001;
			10'd492: USel4 = 4'b0001;
			10'd493: USel4 = 4'b0001;
			10'd494: USel4 = 4'b0001;
			10'd495: USel4 = 4'b0010;
			10'd496: USel4 = 4'b0010;
			10'd497: USel4 = 4'b0010;
			10'd498: USel4 = 4'b0010;
			10'd499: USel4 = 4'b0010;
			10'd500: USel4 = 4'b0010;
			10'd501: USel4 = 4'b0010;
			10'd502: USel4 = 4'b0010;
			10'd503: USel4 = 4'b0010;
			10'd504: USel4 = 4'b0010;
			10'd505: USel4 = 4'b0010;
			10'd506: USel4 = 4'b0000;
			10'd507: USel4 = 4'b0000;
			10'd508: USel4 = 4'b0000;
			10'd509: USel4 = 4'b0000;
			10'd510: USel4 = 4'b0000;
			10'd511: USel4 = 4'b0000;
			10'd512: USel4 = 4'b0000;
			10'd513: USel4 = 4'b0000;
			10'd514: USel4 = 4'b0000;
			10'd515: USel4 = 4'b0000;
			10'd516: USel4 = 4'b0000;
			10'd517: USel4 = 4'b0000;
			10'd518: USel4 = 4'b0100;
			10'd519: USel4 = 4'b0100;
			10'd520: USel4 = 4'b0100;
			10'd521: USel4 = 4'b0100;
			10'd522: USel4 = 4'b0100;
			10'd523: USel4 = 4'b0100;
			10'd524: USel4 = 4'b0100;
			10'd525: USel4 = 4'b0100;
			10'd526: USel4 = 4'b0100;
			10'd527: USel4 = 4'b0100;
			10'd528: USel4 = 4'b0100;
			10'd529: USel4 = 4'b0100;
			10'd530: USel4 = 4'b1000;
			10'd531: USel4 = 4'b1000;
			10'd532: USel4 = 4'b1000;
			10'd533: USel4 = 4'b1000;
			10'd534: USel4 = 4'b1000;
			10'd535: USel4 = 4'b1000;
			10'd536: USel4 = 4'b1000;
			10'd537: USel4 = 4'b1000;
			10'd538: USel4 = 4'b1000;
			10'd539: USel4 = 4'b1000;
			10'd540: USel4 = 4'b1000;
			10'd541: USel4 = 4'b1000;
			10'd542: USel4 = 4'b1000;
			10'd543: USel4 = 4'b1000;
			10'd544: USel4 = 4'b1000;
			10'd545: USel4 = 4'b1000;
			10'd546: USel4 = 4'b1000;
			10'd547: USel4 = 4'b1000;
			10'd548: USel4 = 4'b1000;
			10'd549: USel4 = 4'b1000;
			10'd550: USel4 = 4'b1000;
			10'd551: USel4 = 4'b1000;
			10'd552: USel4 = 4'b1000;
			10'd553: USel4 = 4'b1000;
			10'd554: USel4 = 4'b1000;
			10'd555: USel4 = 4'b1000;
			10'd556: USel4 = 4'b1000;
			10'd557: USel4 = 4'b1000;
			10'd558: USel4 = 4'b1000;
			10'd559: USel4 = 4'b1000;
			10'd560: USel4 = 4'b1000;
			10'd561: USel4 = 4'b1000;
			10'd562: USel4 = 4'b1000;
			10'd563: USel4 = 4'b1000;
			10'd564: USel4 = 4'b1000;
			10'd565: USel4 = 4'b1000;
			10'd566: USel4 = 4'b1000;
			10'd567: USel4 = 4'b1000;
			10'd568: USel4 = 4'b1000;
			10'd569: USel4 = 4'b1000;
			10'd570: USel4 = 4'b1000;
			10'd571: USel4 = 4'b1000;
			10'd572: USel4 = 4'b1000;
			10'd573: USel4 = 4'b1000;
			10'd574: USel4 = 4'b1000;
			10'd575: USel4 = 4'b1000;
			10'd576: USel4 = 4'b0001;
			10'd577: USel4 = 4'b0001;
			10'd578: USel4 = 4'b0001;
			10'd579: USel4 = 4'b0001;
			10'd580: USel4 = 4'b0001;
			10'd581: USel4 = 4'b0001;
			10'd582: USel4 = 4'b0001;
			10'd583: USel4 = 4'b0001;
			10'd584: USel4 = 4'b0001;
			10'd585: USel4 = 4'b0001;
			10'd586: USel4 = 4'b0001;
			10'd587: USel4 = 4'b0001;
			10'd588: USel4 = 4'b0001;
			10'd589: USel4 = 4'b0001;
			10'd590: USel4 = 4'b0001;
			10'd591: USel4 = 4'b0001;
			10'd592: USel4 = 4'b0001;
			10'd593: USel4 = 4'b0001;
			10'd594: USel4 = 4'b0001;
			10'd595: USel4 = 4'b0001;
			10'd596: USel4 = 4'b0001;
			10'd597: USel4 = 4'b0001;
			10'd598: USel4 = 4'b0001;
			10'd599: USel4 = 4'b0001;
			10'd600: USel4 = 4'b0001;
			10'd601: USel4 = 4'b0001;
			10'd602: USel4 = 4'b0001;
			10'd603: USel4 = 4'b0001;
			10'd604: USel4 = 4'b0001;
			10'd605: USel4 = 4'b0001;
			10'd606: USel4 = 4'b0001;
			10'd607: USel4 = 4'b0001;
			10'd608: USel4 = 4'b0001;
			10'd609: USel4 = 4'b0001;
			10'd610: USel4 = 4'b0001;
			10'd611: USel4 = 4'b0001;
			10'd612: USel4 = 4'b0001;
			10'd613: USel4 = 4'b0001;
			10'd614: USel4 = 4'b0001;
			10'd615: USel4 = 4'b0001;
			10'd616: USel4 = 4'b0001;
			10'd617: USel4 = 4'b0001;
			10'd618: USel4 = 4'b0001;
			10'd619: USel4 = 4'b0001;
			10'd620: USel4 = 4'b0001;
			10'd621: USel4 = 4'b0001;
			10'd622: USel4 = 4'b0010;
			10'd623: USel4 = 4'b0010;
			10'd624: USel4 = 4'b0010;
			10'd625: USel4 = 4'b0010;
			10'd626: USel4 = 4'b0010;
			10'd627: USel4 = 4'b0010;
			10'd628: USel4 = 4'b0010;
			10'd629: USel4 = 4'b0010;
			10'd630: USel4 = 4'b0010;
			10'd631: USel4 = 4'b0010;
			10'd632: USel4 = 4'b0010;
			10'd633: USel4 = 4'b0010;
			10'd634: USel4 = 4'b0000;
			10'd635: USel4 = 4'b0000;
			10'd636: USel4 = 4'b0000;
			10'd637: USel4 = 4'b0000;
			10'd638: USel4 = 4'b0000;
			10'd639: USel4 = 4'b0000;
			10'd640: USel4 = 4'b0000;
			10'd641: USel4 = 4'b0000;
			10'd642: USel4 = 4'b0000;
			10'd643: USel4 = 4'b0000;
			10'd644: USel4 = 4'b0000;
			10'd645: USel4 = 4'b0000;
			10'd646: USel4 = 4'b0100;
			10'd647: USel4 = 4'b0100;
			10'd648: USel4 = 4'b0100;
			10'd649: USel4 = 4'b0100;
			10'd650: USel4 = 4'b0100;
			10'd651: USel4 = 4'b0100;
			10'd652: USel4 = 4'b0100;
			10'd653: USel4 = 4'b0100;
			10'd654: USel4 = 4'b0100;
			10'd655: USel4 = 4'b0100;
			10'd656: USel4 = 4'b0100;
			10'd657: USel4 = 4'b0100;
			10'd658: USel4 = 4'b0100;
			10'd659: USel4 = 4'b0100;
			10'd660: USel4 = 4'b1000;
			10'd661: USel4 = 4'b1000;
			10'd662: USel4 = 4'b1000;
			10'd663: USel4 = 4'b1000;
			10'd664: USel4 = 4'b1000;
			10'd665: USel4 = 4'b1000;
			10'd666: USel4 = 4'b1000;
			10'd667: USel4 = 4'b1000;
			10'd668: USel4 = 4'b1000;
			10'd669: USel4 = 4'b1000;
			10'd670: USel4 = 4'b1000;
			10'd671: USel4 = 4'b1000;
			10'd672: USel4 = 4'b1000;
			10'd673: USel4 = 4'b1000;
			10'd674: USel4 = 4'b1000;
			10'd675: USel4 = 4'b1000;
			10'd676: USel4 = 4'b1000;
			10'd677: USel4 = 4'b1000;
			10'd678: USel4 = 4'b1000;
			10'd679: USel4 = 4'b1000;
			10'd680: USel4 = 4'b1000;
			10'd681: USel4 = 4'b1000;
			10'd682: USel4 = 4'b1000;
			10'd683: USel4 = 4'b1000;
			10'd684: USel4 = 4'b1000;
			10'd685: USel4 = 4'b1000;
			10'd686: USel4 = 4'b1000;
			10'd687: USel4 = 4'b1000;
			10'd688: USel4 = 4'b1000;
			10'd689: USel4 = 4'b1000;
			10'd690: USel4 = 4'b1000;
			10'd691: USel4 = 4'b1000;
			10'd692: USel4 = 4'b1000;
			10'd693: USel4 = 4'b1000;
			10'd694: USel4 = 4'b1000;
			10'd695: USel4 = 4'b1000;
			10'd696: USel4 = 4'b1000;
			10'd697: USel4 = 4'b1000;
			10'd698: USel4 = 4'b1000;
			10'd699: USel4 = 4'b1000;
			10'd700: USel4 = 4'b1000;
			10'd701: USel4 = 4'b1000;
			10'd702: USel4 = 4'b1000;
			10'd703: USel4 = 4'b1000;
			10'd704: USel4 = 4'b0001;
			10'd705: USel4 = 4'b0001;
			10'd706: USel4 = 4'b0001;
			10'd707: USel4 = 4'b0001;
			10'd708: USel4 = 4'b0001;
			10'd709: USel4 = 4'b0001;
			10'd710: USel4 = 4'b0001;
			10'd711: USel4 = 4'b0001;
			10'd712: USel4 = 4'b0001;
			10'd713: USel4 = 4'b0001;
			10'd714: USel4 = 4'b0001;
			10'd715: USel4 = 4'b0001;
			10'd716: USel4 = 4'b0001;
			10'd717: USel4 = 4'b0001;
			10'd718: USel4 = 4'b0001;
			10'd719: USel4 = 4'b0001;
			10'd720: USel4 = 4'b0001;
			10'd721: USel4 = 4'b0001;
			10'd722: USel4 = 4'b0001;
			10'd723: USel4 = 4'b0001;
			10'd724: USel4 = 4'b0001;
			10'd725: USel4 = 4'b0001;
			10'd726: USel4 = 4'b0001;
			10'd727: USel4 = 4'b0001;
			10'd728: USel4 = 4'b0001;
			10'd729: USel4 = 4'b0001;
			10'd730: USel4 = 4'b0001;
			10'd731: USel4 = 4'b0001;
			10'd732: USel4 = 4'b0001;
			10'd733: USel4 = 4'b0001;
			10'd734: USel4 = 4'b0001;
			10'd735: USel4 = 4'b0001;
			10'd736: USel4 = 4'b0001;
			10'd737: USel4 = 4'b0001;
			10'd738: USel4 = 4'b0001;
			10'd739: USel4 = 4'b0001;
			10'd740: USel4 = 4'b0001;
			10'd741: USel4 = 4'b0001;
			10'd742: USel4 = 4'b0001;
			10'd743: USel4 = 4'b0001;
			10'd744: USel4 = 4'b0001;
			10'd745: USel4 = 4'b0001;
			10'd746: USel4 = 4'b0001;
			10'd747: USel4 = 4'b0001;
			10'd748: USel4 = 4'b0010;
			10'd749: USel4 = 4'b0010;
			10'd750: USel4 = 4'b0010;
			10'd751: USel4 = 4'b0010;
			10'd752: USel4 = 4'b0010;
			10'd753: USel4 = 4'b0010;
			10'd754: USel4 = 4'b0010;
			10'd755: USel4 = 4'b0010;
			10'd756: USel4 = 4'b0010;
			10'd757: USel4 = 4'b0010;
			10'd758: USel4 = 4'b0010;
			10'd759: USel4 = 4'b0010;
			10'd760: USel4 = 4'b0000;
			10'd761: USel4 = 4'b0000;
			10'd762: USel4 = 4'b0000;
			10'd763: USel4 = 4'b0000;
			10'd764: USel4 = 4'b0000;
			10'd765: USel4 = 4'b0000;
			10'd766: USel4 = 4'b0000;
			10'd767: USel4 = 4'b0000;
			10'd768: USel4 = 4'b0000;
			10'd769: USel4 = 4'b0000;
			10'd770: USel4 = 4'b0000;
			10'd771: USel4 = 4'b0000;
			10'd772: USel4 = 4'b0000;
			10'd773: USel4 = 4'b0000;
			10'd774: USel4 = 4'b0000;
			10'd775: USel4 = 4'b0000;
			10'd776: USel4 = 4'b0100;
			10'd777: USel4 = 4'b0100;
			10'd778: USel4 = 4'b0100;
			10'd779: USel4 = 4'b0100;
			10'd780: USel4 = 4'b0100;
			10'd781: USel4 = 4'b0100;
			10'd782: USel4 = 4'b0100;
			10'd783: USel4 = 4'b0100;
			10'd784: USel4 = 4'b0100;
			10'd785: USel4 = 4'b0100;
			10'd786: USel4 = 4'b0100;
			10'd787: USel4 = 4'b0100;
			10'd788: USel4 = 4'b1000;
			10'd789: USel4 = 4'b1000;
			10'd790: USel4 = 4'b1000;
			10'd791: USel4 = 4'b1000;
			10'd792: USel4 = 4'b1000;
			10'd793: USel4 = 4'b1000;
			10'd794: USel4 = 4'b1000;
			10'd795: USel4 = 4'b1000;
			10'd796: USel4 = 4'b1000;
			10'd797: USel4 = 4'b1000;
			10'd798: USel4 = 4'b1000;
			10'd799: USel4 = 4'b1000;
			10'd800: USel4 = 4'b1000;
			10'd801: USel4 = 4'b1000;
			10'd802: USel4 = 4'b1000;
			10'd803: USel4 = 4'b1000;
			10'd804: USel4 = 4'b1000;
			10'd805: USel4 = 4'b1000;
			10'd806: USel4 = 4'b1000;
			10'd807: USel4 = 4'b1000;
			10'd808: USel4 = 4'b1000;
			10'd809: USel4 = 4'b1000;
			10'd810: USel4 = 4'b1000;
			10'd811: USel4 = 4'b1000;
			10'd812: USel4 = 4'b1000;
			10'd813: USel4 = 4'b1000;
			10'd814: USel4 = 4'b1000;
			10'd815: USel4 = 4'b1000;
			10'd816: USel4 = 4'b1000;
			10'd817: USel4 = 4'b1000;
			10'd818: USel4 = 4'b1000;
			10'd819: USel4 = 4'b1000;
			10'd820: USel4 = 4'b1000;
			10'd821: USel4 = 4'b1000;
			10'd822: USel4 = 4'b1000;
			10'd823: USel4 = 4'b1000;
			10'd824: USel4 = 4'b1000;
			10'd825: USel4 = 4'b1000;
			10'd826: USel4 = 4'b1000;
			10'd827: USel4 = 4'b1000;
			10'd828: USel4 = 4'b1000;
			10'd829: USel4 = 4'b1000;
			10'd830: USel4 = 4'b1000;
			10'd831: USel4 = 4'b1000;
			10'd832: USel4 = 4'b0001;
			10'd833: USel4 = 4'b0001;
			10'd834: USel4 = 4'b0001;
			10'd835: USel4 = 4'b0001;
			10'd836: USel4 = 4'b0001;
			10'd837: USel4 = 4'b0001;
			10'd838: USel4 = 4'b0001;
			10'd839: USel4 = 4'b0001;
			10'd840: USel4 = 4'b0001;
			10'd841: USel4 = 4'b0001;
			10'd842: USel4 = 4'b0001;
			10'd843: USel4 = 4'b0001;
			10'd844: USel4 = 4'b0001;
			10'd845: USel4 = 4'b0001;
			10'd846: USel4 = 4'b0001;
			10'd847: USel4 = 4'b0001;
			10'd848: USel4 = 4'b0001;
			10'd849: USel4 = 4'b0001;
			10'd850: USel4 = 4'b0001;
			10'd851: USel4 = 4'b0001;
			10'd852: USel4 = 4'b0001;
			10'd853: USel4 = 4'b0001;
			10'd854: USel4 = 4'b0001;
			10'd855: USel4 = 4'b0001;
			10'd856: USel4 = 4'b0001;
			10'd857: USel4 = 4'b0001;
			10'd858: USel4 = 4'b0001;
			10'd859: USel4 = 4'b0001;
			10'd860: USel4 = 4'b0001;
			10'd861: USel4 = 4'b0001;
			10'd862: USel4 = 4'b0001;
			10'd863: USel4 = 4'b0001;
			10'd864: USel4 = 4'b0001;
			10'd865: USel4 = 4'b0001;
			10'd866: USel4 = 4'b0001;
			10'd867: USel4 = 4'b0001;
			10'd868: USel4 = 4'b0001;
			10'd869: USel4 = 4'b0001;
			10'd870: USel4 = 4'b0001;
			10'd871: USel4 = 4'b0001;
			10'd872: USel4 = 4'b0001;
			10'd873: USel4 = 4'b0001;
			10'd874: USel4 = 4'b0010;
			10'd875: USel4 = 4'b0010;
			10'd876: USel4 = 4'b0010;
			10'd877: USel4 = 4'b0010;
			10'd878: USel4 = 4'b0010;
			10'd879: USel4 = 4'b0010;
			10'd880: USel4 = 4'b0010;
			10'd881: USel4 = 4'b0010;
			10'd882: USel4 = 4'b0010;
			10'd883: USel4 = 4'b0010;
			10'd884: USel4 = 4'b0010;
			10'd885: USel4 = 4'b0010;
			10'd886: USel4 = 4'b0010;
			10'd887: USel4 = 4'b0010;
			10'd888: USel4 = 4'b0000;
			10'd889: USel4 = 4'b0000;
			10'd890: USel4 = 4'b0000;
			10'd891: USel4 = 4'b0000;
			10'd892: USel4 = 4'b0000;
			10'd893: USel4 = 4'b0000;
			10'd894: USel4 = 4'b0000;
			10'd895: USel4 = 4'b0000;
			10'd896: USel4 = 4'b0000;
			10'd897: USel4 = 4'b0000;
			10'd898: USel4 = 4'b0000;
			10'd899: USel4 = 4'b0000;
			10'd900: USel4 = 4'b0000;
			10'd901: USel4 = 4'b0000;
			10'd902: USel4 = 4'b0000;
			10'd903: USel4 = 4'b0000;
			10'd904: USel4 = 4'b0100;
			10'd905: USel4 = 4'b0100;
			10'd906: USel4 = 4'b0100;
			10'd907: USel4 = 4'b0100;
			10'd908: USel4 = 4'b0100;
			10'd909: USel4 = 4'b0100;
			10'd910: USel4 = 4'b0100;
			10'd911: USel4 = 4'b0100;
			10'd912: USel4 = 4'b0100;
			10'd913: USel4 = 4'b0100;
			10'd914: USel4 = 4'b0100;
			10'd915: USel4 = 4'b0100;
			10'd916: USel4 = 4'b0100;
			10'd917: USel4 = 4'b0100;
			10'd918: USel4 = 4'b0100;
			10'd919: USel4 = 4'b0100;
			10'd920: USel4 = 4'b1000;
			10'd921: USel4 = 4'b1000;
			10'd922: USel4 = 4'b1000;
			10'd923: USel4 = 4'b1000;
			10'd924: USel4 = 4'b1000;
			10'd925: USel4 = 4'b1000;
			10'd926: USel4 = 4'b1000;
			10'd927: USel4 = 4'b1000;
			10'd928: USel4 = 4'b1000;
			10'd929: USel4 = 4'b1000;
			10'd930: USel4 = 4'b1000;
			10'd931: USel4 = 4'b1000;
			10'd932: USel4 = 4'b1000;
			10'd933: USel4 = 4'b1000;
			10'd934: USel4 = 4'b1000;
			10'd935: USel4 = 4'b1000;
			10'd936: USel4 = 4'b1000;
			10'd937: USel4 = 4'b1000;
			10'd938: USel4 = 4'b1000;
			10'd939: USel4 = 4'b1000;
			10'd940: USel4 = 4'b1000;
			10'd941: USel4 = 4'b1000;
			10'd942: USel4 = 4'b1000;
			10'd943: USel4 = 4'b1000;
			10'd944: USel4 = 4'b1000;
			10'd945: USel4 = 4'b1000;
			10'd946: USel4 = 4'b1000;
			10'd947: USel4 = 4'b1000;
			10'd948: USel4 = 4'b1000;
			10'd949: USel4 = 4'b1000;
			10'd950: USel4 = 4'b1000;
			10'd951: USel4 = 4'b1000;
			10'd952: USel4 = 4'b1000;
			10'd953: USel4 = 4'b1000;
			10'd954: USel4 = 4'b1000;
			10'd955: USel4 = 4'b1000;
			10'd956: USel4 = 4'b1000;
			10'd957: USel4 = 4'b1000;
			10'd958: USel4 = 4'b1000;
			10'd959: USel4 = 4'b1000;
			10'd960: USel4 = 4'b0001;
			10'd961: USel4 = 4'b0001;
			10'd962: USel4 = 4'b0001;
			10'd963: USel4 = 4'b0001;
			10'd964: USel4 = 4'b0001;
			10'd965: USel4 = 4'b0001;
			10'd966: USel4 = 4'b0001;
			10'd967: USel4 = 4'b0001;
			10'd968: USel4 = 4'b0001;
			10'd969: USel4 = 4'b0001;
			10'd970: USel4 = 4'b0001;
			10'd971: USel4 = 4'b0001;
			10'd972: USel4 = 4'b0001;
			10'd973: USel4 = 4'b0001;
			10'd974: USel4 = 4'b0001;
			10'd975: USel4 = 4'b0001;
			10'd976: USel4 = 4'b0001;
			10'd977: USel4 = 4'b0001;
			10'd978: USel4 = 4'b0001;
			10'd979: USel4 = 4'b0001;
			10'd980: USel4 = 4'b0001;
			10'd981: USel4 = 4'b0001;
			10'd982: USel4 = 4'b0001;
			10'd983: USel4 = 4'b0001;
			10'd984: USel4 = 4'b0001;
			10'd985: USel4 = 4'b0001;
			10'd986: USel4 = 4'b0001;
			10'd987: USel4 = 4'b0001;
			10'd988: USel4 = 4'b0001;
			10'd989: USel4 = 4'b0001;
			10'd990: USel4 = 4'b0001;
			10'd991: USel4 = 4'b0001;
			10'd992: USel4 = 4'b0001;
			10'd993: USel4 = 4'b0001;
			10'd994: USel4 = 4'b0001;
			10'd995: USel4 = 4'b0001;
			10'd996: USel4 = 4'b0001;
			10'd997: USel4 = 4'b0001;
			10'd998: USel4 = 4'b0001;
			10'd999: USel4 = 4'b0001;
			10'd1000: USel4 = 4'b0001;
			10'd1001: USel4 = 4'b0001;
			10'd1002: USel4 = 4'b0010;
			10'd1003: USel4 = 4'b0010;
			10'd1004: USel4 = 4'b0010;
			10'd1005: USel4 = 4'b0010;
			10'd1006: USel4 = 4'b0010;
			10'd1007: USel4 = 4'b0010;
			10'd1008: USel4 = 4'b0010;
			10'd1009: USel4 = 4'b0010;
			10'd1010: USel4 = 4'b0010;
			10'd1011: USel4 = 4'b0010;
			10'd1012: USel4 = 4'b0010;
			10'd1013: USel4 = 4'b0010;
			10'd1014: USel4 = 4'b0010;
			10'd1015: USel4 = 4'b0010;
			10'd1016: USel4 = 4'b0000;
			10'd1017: USel4 = 4'b0000;
			10'd1018: USel4 = 4'b0000;
			10'd1019: USel4 = 4'b0000;
			10'd1020: USel4 = 4'b0000;
			10'd1021: USel4 = 4'b0000;
			10'd1022: USel4 = 4'b0000;
			10'd1023: USel4 = 4'b0000;
		endcase
	end
	always @(*) begin
		if (_sv2v_0)
			;
		if (Sqrt) begin
			if (j1)
				A = 3'b101;
			else if (Smsbs[4] == 1)
				A = 3'b111;
			else
				A = Smsbs[2:0];
		end
		else
			A = Dmsbs;
	end
	assign udigit = (Sqrt & j0 ? 4'b0100 : USel4);
	initial _sv2v_0 = 0;
endmodule
